//==================================================================================================
//  Filename      : tb_FPU_PIPELINED_FPADDSUB2_vector_testing.v
//  Created On    : 2016-09-24 01:24:56
//  Last Modified : 2016-09-24 01:24:56
//  Revision      :
//  Author        : Jorge Sequeira Rojas
//  Company       : Instituto Tecnologico de Costa Rica
//  Email         : jsequeira@gmail.com
//
//  Description   :
//
//
//==================================================================================================

`timescale 1ns/1ps


module tb_FPU_PIPELINED_FPADDSUB2_vector_testing (); /* this is automatically generated */

  localparam PERIOD = 10;

  // (*NOTE*) replace reset, clock
   parameter W = 32;
   parameter EW = 8;
   parameter SW = 23;
   parameter SWR=26;
   parameter EWR = 5;  //Single Precision */

  // parameter W   = 64;
  // parameter EW  = 11;
  // parameter SW  = 52;
  // parameter SWR = 55;
  // parameter EWR = 6;

  reg         clk;
  reg         rst;
  reg         beg_OP;
  reg [W-1:0] Data_X;
  reg [W-1:0] Data_Y;
  reg         add_subt;
  wire        busy;
  wire        overflow_flag;
  wire        underflow_flag;
  wire        zero_flag;

  wire [W-1:0] final_result_ieee;
  reg [SW-1:0] final_result_ieee_mantissa;
  reg [EW-1:0] final_result_ieee_exponent;
  reg          final_result_ieee_sign;

  wire ready;

//Temps for the testbench and verification

  reg [SW-1:0] Data_X_mant;
  reg [SW-1:0] Data_Y_mant;
  reg [EW-1:0] Data_X_exp;
  reg [EW-1:0] Data_Y_exp;
  reg Data_X_sign;
  reg Data_Y_sign;

  reg  [W-1:0] formatted_number_W;
  reg overflow_flag_t, underflow_flag_t;

  reg [EWR-1:0] LZD_raw_val_EWR;
  reg [W-1:0]  Theoretical_result;
  reg [SW-1:0] Theoretical_result_mantissa;
  reg [EW-1:0] Theoretical_result_exponent;
  reg Theoretical_result_sign;

  reg [W-1:0] Array_IN [0:((2**PERIOD)-1)];
  reg [W-1:0] Array_IN_2 [0:((2**PERIOD)-1)];
  integer contador;
  integer FileSaveData;
  integer Cont_CLK;
  integer Recept;

  FPU_PIPELINED_FPADDSUB #(
      .W(W),
      .EW(EW),
      .SW(SW),
      .SWR(SWR),
      .EWR(EWR)
    ) inst_FPU_PIPELINED_FPADDSUB (
      .clk               (clk),
      .rst               (rst),
      .beg_OP            (beg_OP),
      .Data_X            (Data_X),
      .Data_Y            (Data_Y),
      .add_subt          (add_subt),
      .busy              (busy),
      .overflow_flag     (overflow_flag),
      .underflow_flag    (underflow_flag),
      .zero_flag         (zero_flag),
      .ready             (ready),
      .final_result_ieee (final_result_ieee)
    );

always begin
    #1;
    final_result_ieee_mantissa = final_result_ieee[SW-1:0];
    final_result_ieee_exponent = final_result_ieee[W-2:SW];
    final_result_ieee_sign     = final_result_ieee[W-1];
    Data_X_mant = Data_X[SW-1:0];
    Data_Y_mant = Data_Y[SW-1:0];
    Data_X_exp  = Data_X[W-2:SW];
    Data_Y_exp  = Data_Y[W-2:SW];
    Data_X_sign = Data_X[W-1];
    Data_Y_sign = Data_Y[W-1];
    Theoretical_result_mantissa = Theoretical_result[SW-1:0];
    Theoretical_result_exponent = Theoretical_result[W-2:SW];
    Theoretical_result_sign = Theoretical_result[W-1];

end

// function [EWR-1:0] LZD_raw; // function definition starts here
//    input [SWR-1:0] ADD_SUB_RAW;
//    integer k;
//    begin
//      LZD_raw = 0;
//      k=SWR-1;
//      while(ADD_SUB_RAW[k] == 0) begin
//        k = k-1;
//        LZD_raw = LZD_raw + 1;
//         $display("This is the bit analized %d", k);
//         $display("This is the bit analized %d", ADD_SUB_RAW[k]);
//         $display("Number of 0s %d", LZD_raw);
//      end
//    end
//  endfunction


   initial begin
    FileSaveData = $fopen("ResultadoXilinxFLM.txt","w");
    rst = 1;
    add_subt = 0;
    beg_OP = 0;
    Data_Y = 0;
    Data_X = 0;
    Data_X_mant = 0;
    Data_Y_mant = 0;
    Data_X_exp  = 0;
    Data_Y_exp  = 0;
    Data_X_sign = 0;
    Data_Y_sign = 0;
    Theoretical_result = 32'hbe1abef8;
    //Inicializa las variables del testbench
    contador = 0;
    Cont_CLK = 0;
    Recept = 1;


    #100 rst = 0;


   end

   //**************************** Se lee el archivo txt y se almacena en un arrays***************************************************//

    initial begin
        $readmemh("Hexadecimal_A.txt", Array_IN);
        $readmemh("Hexadecimal_B.txt", Array_IN_2);
    end

     //**************************** Transmision de datos de forma paralela ************************************************************//

  always @(negedge clk) begin
      if (contador == (2**PERIOD)) begin
          $fclose(FileSaveData);
          $finish;
      end else if(ready) begin
        $fwrite(FileSaveData,"%h\n",final_result_ieee);
      end

  end

always @(negedge clk) begin
    if(rst) begin
        contador = 0;
    end
    else if(~busy) begin
        Data_X = Array_IN[contador];
        Data_Y = Array_IN_2[contador];
        contador = contador + 1;
        beg_OP = 1;
    end
end

  // clock

  initial begin
    clk = 0;
    forever #(PERIOD/2) clk = ~clk;
  end

endmodule


